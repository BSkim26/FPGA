`timescale 1ns / 1ps

module tb_Microprocessor();                                         //TEST Bench
    reg clk,clk_10;                                                 //�Է°� ��� ����
    reg [3:0] sw;    
    reg [3:0] btn;         
    wire [3:0] led;           
    wire [1:0] seg_en;       
    wire [6:0] seg_ab, seg_cd;

Microprocessor uut(clk,clk_10,sw,btn,led,seg_en,seg_ab,seg_cd);     //Microprocessor module ����

always #5 clk = ~clk;                                               // 100MHz�� clk ����
always #50 clk_10 = ~clk_10;                                        // Overflow�� ���� 10Hz clk ����


initial begin
    clk=0;clk_10=0;btn=0;sw=0;                                      // �ʱⰪ ����
    
    #100                                                            // implementation �ʱ� delay ������ 100ns delay 
    #10                   btn[0] = 1'b1;                            // ADDI $1, 5, $1(1100_0001_0101_0001)
    #10                   btn[0] = 1'b0;  
    #10     sw = 4'b1100;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0001;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0101;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0001;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0000;
    #10
    #50                    btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10
    #10
    
    #10                    btn[0] = 1'b1;                           // SUBI $2, 6, $2(1101_0010_0110_0010)
    #10                   btn[0] = 1'b0;  
    #10     sw = 4'b1101;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0010;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0110;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0010;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0000;
    #10
    #50                    btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10
    #10
    
    #10                    btn[0] = 1'b1;                           // ADD $1, $2, $3(1010_0001_0010_0011)
    #10                   btn[0] = 1'b0;  
    #10     sw = 4'b1010;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0001;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0010;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0011;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0000;
    #10
    #50                    btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10
    #10
    
    #10                    btn[0] = 1'b1;                           // NOP x x x(0000_xxxx_xxxx_xxxx)
    #10                   btn[0] = 1'b0;  
    #10     sw = 4'b0000;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0001;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0010;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0011;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0000;
    #10
    #50                    btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10
    #10
    
    #10                    btn[0] = 1'b1;                           // Write  x, 7, $4(0001_xxxx_0111_0100)
    #10                   btn[0] = 1'b0;  
    #10     sw = 4'b0001;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0001;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0111;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0100;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0000;
    #10
    #50                    btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10
    #10
    
    #10                    btn[0] = 1'b1;                           // SUB $4, $2, $5(1011_0100_0010_0101)
    #10                   btn[0] = 1'b0;  
    #10     sw = 4'b1011;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0100;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0010;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0101;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0000;
    #10
    #610                    btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10
    #10

    #10                    btn[0] = 1'b1;                           // NOT $3, x, $5(0100_0011_xxxx_0101)
    #10                   btn[0] = 1'b0;  
    #10     sw = 4'b0100;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0011;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0111;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0101;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0000;
    #10
    #50                    btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10
    #10
    
    #10                    btn[0] = 1'b1;                           // XOR $1, $3, $1(0111_0001_0011_0001)
    #10                   btn[0] = 1'b0;  
    #10     sw = 4'b0111;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0001;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0011;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0001;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0000;
    #10
    #50                    btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10
    #10
    
    #10                    btn[0] = 1'b1;                           // NOR $2, $5, $5(1001_0010_0101_0101)
    #10                   btn[0] = 1'b0;  
    #10     sw = 4'b1001;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0010;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0101;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0101;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0000;
    #10
    #50                    btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10
    #10
    
    #10                    btn[0] = 1'b1;                           // Read $2, x, x(0010_0010_xxxx_xxxx)
    #10                   btn[0] = 1'b0;  
    #10     sw = 4'b0010;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0010;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b1110;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0100;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0000;
    #10
    #50                    btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10
    #10
    
    #10                    btn[0] = 1'b1;                           // NAND $3, $1, $2(1000_0011_0001_0010)
    #10                   btn[0] = 1'b0;  
    #10     sw = 4'b1000;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0011;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0001;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0010;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0000;
    #10
    #50                    btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10
    #10
    
    #10                    btn[0] = 1'b1;                           // Left Shift $2, 3, $0(1110_0010_0011_0000)
    #10                   btn[0] = 1'b0;  
    #10     sw = 4'b1110;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0010;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0011;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0000;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0000;
    #10
    #50                    btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10
    #10
    
    #10                    btn[0] = 1'b1;                           // Copy $3, x, $4(0011_0011_xxxx_0100)
    #10                   btn[0] = 1'b0;  
    #10     sw = 4'b0011;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0011;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b1010;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0100;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0000;
    #10
    #50                    btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10
    #10
    
    #10                    btn[0] = 1'b1;                           // AND $1, $2, $3(0101_0001_0010_0011)
    #10                   btn[0] = 1'b0;  
    #10     sw = 4'b0101;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0001;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0010;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0011;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0000;
    #10
    #50                    btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10
    #10
    
    #10                    btn[0] = 1'b1;                           // ADD $2, $2, $2(1010_0010_0010_0010)
    #10                   btn[0] = 1'b0;  
    #10     sw = 4'b1010;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0010;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0010;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0010;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0000;
    #10
    #610                    btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10
    #10
    
    #10                    btn[0] = 1'b1;                           // OR $2, $1, $1(0110_0010_0001_0001)
    #10                   btn[0] = 1'b0;  
    #10     sw = 4'b0110;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0010;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0001;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0001;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0000;
    #10
    #50                    btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10
    #10
    
    #10                    btn[0] = 1'b1;                           // Shift Right $2, 1, $5(1111_0010_0001_0101)
    #10                   btn[0] = 1'b0;  
    #10     sw = 4'b1111;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0010;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0001;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0101;  btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10     sw = 4'b0000;
    #10
    #50                    btn[0] = 1'b1;
    #10                   btn[0] = 1'b0;
    #10
    #10;
end

endmodule
