`timescale 1ns / 1ps



module MUX8bit(
    input [7:0] a,      // 8bit�� �Է��� �ޱ� ���� 8bit a�� input���� �����Ѵ�.
    input [2:0] sel,    // �Է��� ������ ����� �� �ֵ��� 3bit sel�� �����Ѵ�.
    output  out         // out�� output �������� �����Ѵ�.
    );
    
    assign out =    (sel==3'b000) ? a[0] :          // sel�� 000�̶�� a[0]�� ����Ѵ�.
                    (sel==3'b001) ? a[1] :          // sel�� 001�̶�� a[1]�� ����Ѵ�.
                    (sel==3'b010) ? a[2] :          // sel�� 010�̶�� a[2]�� ����Ѵ�.
                    (sel==3'b011) ? a[3] :          // sel�� 011�̶�� a[3]�� ����Ѵ�.
                    (sel==3'b100) ? a[4] :          //sel�� 100�̶�� a[4]�� ����Ѵ�.
                    (sel==3'b101) ? a[5] :          //sel�� 000�̶�� a[5]�� ����Ѵ�.
                    (sel==3'b110) ? a[6] :          //sel�� 110�̶�� a[6]�� ����Ѵ�.
                    (sel==3'b111) ? a[7] : 1'bx;    //sel�� 111�̶�� a[7]�� ����ϰ� �� �̿��� ���� �ԷµǸ� x�� ����Ѵ�.
endmodule